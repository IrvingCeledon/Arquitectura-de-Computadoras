// 1.- Module definition - inputs and outputs.
module _and (input A, input B, output C);
  
// 2.- Signals and internal elements.
// N/A
  
// 3.- Module behavior
//     (assignments, instances, connections, etc).
assign  C = A&B;

endmodule
