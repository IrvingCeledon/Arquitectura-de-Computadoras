module Burrito (DIR
