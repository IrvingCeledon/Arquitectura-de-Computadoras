// 1.- Module definition - input and output

module _and (input A, input B, output C);
// 2.- Signals and intern elements
// N/A
// 3.- Module behaviour
//     (assignaments, instances, connections, etc).

assign  C = A&B;

endmodule